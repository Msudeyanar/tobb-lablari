module moduleName (        
        input A,
        input B,
        input Cin,
        output S,

        output Cout, 

)


   




endmodule
